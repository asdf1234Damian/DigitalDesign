module converter ( 
	i,
	c,
	o
	) ;

input [8:0] i;
input  c;
inout [8:0] o;
