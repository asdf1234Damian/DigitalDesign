module converter ( 
	i,
	c,
	o
	) ;

input [7:0] i;
input  c;
inout [7:0] o;
