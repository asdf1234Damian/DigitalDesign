module holapalabra ( 
	invec,
	control,
	outvec
	) ;

input [3:0] invec;
input  control;
inout [6:0] outvec;
