module encoder ( 
	i,
	o
	) ;

input [9:0] i;
inout [3:0] o;
