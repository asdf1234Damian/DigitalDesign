module fft ( 
	toggle,
	clr,
	pre,
	clock,
	q,
	nq
	) ;

input  toggle;
input  clr;
input  pre;
input  clock;
inout  q;
inout  nq;
