module encoder ( 
	input,
	output
	) ;

input [9:0] input;
inout [3:0] output;
