module decoder ( 
	i,
	c,
	o
	) ;

input [3:0] i;
input  c;
inout [6:0] o;
