module converter ( 
	i,
	c,
	o
	) ;

input [3:0] i;
input  c;
inout [3:0] o;
