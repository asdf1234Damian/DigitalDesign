library ieee;
use ieee.std_logic_1164.all;

entity seisEntradas is
  port (
  a,b,c,d,e,f: in std_logic;
  z: out std_logic
  );
end entity;

