architecture XorOperaciones of SeisEntradas is 
begin 
z<=((((a xor b) xor c)xor d)xor e)xor f;
end architecture;